library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity transfer is
	generic(
		framlent:integer:=8
	);
	Port(
		bclkt				: in std_logic;
		resett				: in std_logic;
		xmit_cmd_p			: in std_logic;
		buf0				: in std_logic_vector(7 downto 0);
        buf1				: in std_logic_vector(7 downto 0);
        buf2				: in std_logic_vector(7 downto 0);
        buf3				: in std_logic_vector(7 downto 0);
        buf4				: in std_logic_vector(7 downto 0);
		txd					: out std_logic;
		txd_done			: out std_logic 
	);
end transfer;

architecture behave of transfer is
	type states is (x_idle,x_start,x_wait,x_shift,x_stop);                --??????????
	signal state	: states := x_idle;

begin
	process(bclkt, resett, xmit_cmd_p)                         --????????????????
		variable xcnt16		: std_logic_vector(4 downto 0) 	:= "00000";            --?????��?????
		variable xbitcnt	: integer:=0;
		variable txds		: std_logic;
		variable buf		: std_logic_vector(7 downto 0);
        variable cnt        : integer := 0;
	begin
		if resett='0' then
			state <= x_idle;
			txd_done <= '1';
			txds := '1';           --??��
			cnt := 0;
		elsif rising_edge(bclkt) then
			case state is
				when x_idle =>	--??1??????????????????
					txd_done <= '1';
					if xmit_cmd_p='1' then
						state <= x_start;
						txd_done <= '0';
					else
						state <= x_idle;
					end if;
				when x_start =>	--??2??????????????��
                    case cnt is
                        when 0 => buf := buf0;
                        when 1 => buf := buf1;
                        when 2 => buf := buf2;
                        when 3 => buf := buf3;
                        when 4 => buf := buf4;
                        when others => buf := buf0;
                    end case;
					state <= x_wait;
					xcnt16 := "00000";
					txds := '0';
				when x_wait =>	--??3???????
					if xcnt16 >= "01110" then
						if xbitcnt=framlent then
							state <= x_stop;
							xbitcnt := 0;
						else
							state <= x_shift;
						end if;
						xcnt16 := "00000";
					else
						xcnt16 := xcnt16+1;
						state <= x_wait;
					end if;
				when x_shift =>
					txds := buf(xbitcnt);
					xbitcnt := xbitcnt+1;
					state <= x_wait;				                                        --??4??????????????��??????
				when x_stop =>                         --??5????��??????
					if xcnt16 >= "01111" then
                        if cnt < 4 then
                            cnt := cnt + 1;
                            xcnt16 := "00000";
                            state <= x_start;
                        else
                            txd_done <= '1';
                            if xmit_cmd_p = '0' then
                                cnt := 0;
                                state <= x_idle;
                            else
    							xcnt16 := xcnt16;
    							state <= x_stop;
                            end if;
                        end if;
					else
						xcnt16 := xcnt16+1;
						txds := '1';
						state <= x_stop;
					end if;
				when others =>
					state <= x_idle;
			end case;
		end if;
		txd <= txds;
	end process;
end behave;
