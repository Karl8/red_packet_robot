library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package definitions is
    constant data_width : integer := 8; 
    constant address_width : integer := 16;
end package definitions;
